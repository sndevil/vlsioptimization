module F291 (b , e , VV291V); 
input b , e;
output VV291V;
and f0 (VV291V , b , e);
endmodule