module F117 (a , b , VV117V); 
input a , b;
output VV117V;
or f0 (VV117V , a , b);
endmodule