module F201 (VV197V , VV200V , VV201V); 
input VV197V , VV200V;
output VV201V;
xor f0 (VV201V , VV197V , VV200V);
endmodule