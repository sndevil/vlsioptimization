module F364 (b , e , VV364V); 
input b , e;
output VV364V;
xor f0 (VV364V , b , e);
endmodule