module F227 (b , d , VV227V); 
input b , d;
output VV227V;
and f0 (VV227V , b , d);
endmodule