module F49 (VV47V , VV48V , VV49V); 
input VV47V , VV48V;
output VV49V;
and f0 (VV49V , VV47V , VV48V);
endmodule