module F20 (b , d , VV20V); 
input b , d;
output VV20V;
or f0 (VV20V , b , d);
endmodule