module F65 (d , c , VV65V); 
input d , c;
output VV65V;
wire WW64W0W;

not f0 (WW64W0W , d);
and f1 (VV65V , WW64W0W , c);
endmodule