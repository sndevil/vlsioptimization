module F143 (e , a , VV143V); 
input e , a;
output VV143V;
xor f0 (VV143V , e , a);
endmodule