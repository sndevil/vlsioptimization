module F23 (c , e , VV23V); 
input c , e;
output VV23V;
xor f0 (VV23V , c , e);
endmodule