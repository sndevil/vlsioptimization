module F114 (d , a , VV114V); 
input d , a;
output VV114V;
xor f0 (VV114V , d , a);
endmodule