module F32 (e , c , VV32V); 
input e , c;
output VV32V;
or f0 (VV32V , e , c);
endmodule