module F5 (e , k , VV5V); 
input e , k;
output VV5V;
xor f0 (VV5V , e , k);
endmodule