module F121 (a , c , VV121V); 
input a , c;
output VV121V;
or f0 (VV121V , a , c);
endmodule