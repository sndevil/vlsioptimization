module F99 (c , d , VV99V); 
input c , d;
output VV99V;
or f0 (VV99V , c , d);
endmodule