module F171 (VV163V , VV170V , VV171V); 
input VV163V , VV170V;
output VV171V;
or f0 (VV171V , VV163V , VV170V);
endmodule