module F5 (a , b , VV5V); 
input a , b;
output VV5V;
xor f0 (VV5V , a , b);
endmodule