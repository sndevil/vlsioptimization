module F48 (b , c , VV48V); 
input b , c;
output VV48V;
and f0 (VV48V , b , c);
endmodule