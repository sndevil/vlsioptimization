module F14 (VV10V , VV13V , VV14V); 
input VV10V , VV13V;
output VV14V;
and f0 (VV14V , VV10V , VV13V);
endmodule