module F216 (a , c , VV216V); 
input a , c;
output VV216V;
and f0 (VV216V , a , c);
endmodule