module F76 (VV74V , VV75V , VV76V); 
input VV74V , VV75V;
output VV76V;
or f0 (VV76V , VV74V , VV75V);
endmodule