module F136 (d , e , VV136V); 
input d , e;
output VV136V;
and f0 (VV136V , d , e);
endmodule