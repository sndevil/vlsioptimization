module F138 (c , d , VV138V); 
input c , d;
output VV138V;
xor f0 (VV138V , c , d);
endmodule