module F1 (d , r , VV1V); 
input d , r;
output VV1V;
and f0 (VV1V , d , r);
endmodule