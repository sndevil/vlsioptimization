module F70 (d , c , VV70V); 
input d , c;
output VV70V;
wire WW69W0W;

not f0 (WW69W0W , d);
or f1 (VV70V , WW69W0W , c);
endmodule