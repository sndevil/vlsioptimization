module F73 (c , a , VV73V); 
input c , a;
output VV73V;
xor f0 (VV73V , c , a);
endmodule