module F361 (VV353V , VV360V , VV361V); 
input VV353V , VV360V;
output VV361V;
xor f0 (VV361V , VV353V , VV360V);
endmodule