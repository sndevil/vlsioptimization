module F77 (VV75V , VV76V , VV77V); 
input VV75V , VV76V;
output VV77V;
and f0 (VV77V , VV75V , VV76V);
endmodule