module F151 (d , b , VV151V); 
input d , b;
output VV151V;
or f0 (VV151V , d , b);
endmodule