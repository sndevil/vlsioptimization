module F51 (e , b , VV51V); 
input e , b;
output VV51V;
or f0 (VV51V , e , b);
endmodule