module F62 (a , c , VV62V); 
input a , c;
output VV62V;
and f0 (VV62V , a , c);
endmodule