module F166 (VV164V , VV165V , VV166V); 
input VV164V , VV165V;
output VV166V;
xor f0 (VV166V , VV164V , VV165V);
endmodule