module F9 (c , d , VV9V); 
input c , d;
output VV9V;
xor f0 (VV9V , c , d);
endmodule