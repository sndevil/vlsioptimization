module F71 (VV69V , VV70V , VV71V); 
input VV69V , VV70V;
output VV71V;
xor f0 (VV71V , VV69V , VV70V);
endmodule