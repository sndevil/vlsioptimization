module F246 (d , c , VV246V); 
input d , c;
output VV246V;
xor f0 (VV246V , d , c);
endmodule