module F55 (a , e , VV55V); 
input a , e;
output VV55V;
or f0 (VV55V , a , e);
endmodule