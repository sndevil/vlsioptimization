module F33 (VV31V , VV32V , VV33V); 
input VV31V , VV32V;
output VV33V;
or f0 (VV33V , VV31V , VV32V);
endmodule