module F162 (VV160V , VV161V , VV162V); 
input VV160V , VV161V;
output VV162V;
and f0 (VV162V , VV160V , VV161V);
endmodule