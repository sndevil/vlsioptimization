module F259 (a , b , VV259V); 
input a , b;
output VV259V;
and f0 (VV259V , a , b);
endmodule