module F99 (VV97V , VV98V , VV99V); 
input VV97V , VV98V;
output VV99V;
or f0 (VV99V , VV97V , VV98V);
endmodule