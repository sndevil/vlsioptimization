module F186 (VV182V , VV185V , VV186V); 
input VV182V , VV185V;
output VV186V;
or f0 (VV186V , VV182V , VV185V);
endmodule