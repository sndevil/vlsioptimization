module F19 (c , e , VV19V); 
input c , e;
output VV19V;
or f0 (VV19V , c , e);
endmodule