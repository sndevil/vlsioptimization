module F172 (VV156V' , VV171V , VV172V); 
input VV156V' , VV171V;
output VV172V;
and f0 (VV172V , VV156V' , VV171V);
endmodule