module F4 (f , n , VV4V); 
input f , n;
output VV4V;
or f0 (VV4V , f , n);
endmodule