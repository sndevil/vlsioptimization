module F104 (a , e , VV104V); 
input a , e;
output VV104V;
and f0 (VV104V , a , e);
endmodule