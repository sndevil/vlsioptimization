module F392 (VV384V , VV391V , VV392V); 
input VV384V , VV391V;
output VV392V;
or f0 (VV392V , VV384V , VV391V);
endmodule