module F195 (VV187V , VV194V , VV195V); 
input VV187V , VV194V;
output VV195V;
or f0 (VV195V , VV187V , VV194V);
endmodule