module F393 (VV377V , VV392V , VV393V); 
input VV377V , VV392V;
output VV393V;
or f0 (VV393V , VV377V , VV392V);
endmodule