module F100 (VV98V , VV99V , VV100V); 
input VV98V , VV99V;
output VV100V;
or f0 (VV100V , VV98V , VV99V);
endmodule