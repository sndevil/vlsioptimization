module F109 (VV101V , VV108V , VV109V); 
input VV101V , VV108V;
output VV109V;
or f0 (VV109V , VV101V , VV108V);
endmodule