module F36 (VV34V , VV35V , VV36V); 
input VV34V , VV35V;
output VV36V;
xor f0 (VV36V , VV34V , VV35V);
endmodule