module F374 (e , d , VV374V); 
input e , d;
output VV374V;
and f0 (VV374V , e , d);
endmodule