module F103 (c , d , VV103V); 
input c , d;
output VV103V;
and f0 (VV103V , c , d);
endmodule