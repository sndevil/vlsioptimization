module F214 (VV212V , VV213V , VV214V); 
input VV212V , VV213V;
output VV214V;
or f0 (VV214V , VV212V , VV213V);
endmodule