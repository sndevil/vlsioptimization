module F27 (d , c , VV27V); 
input d , c;
output VV27V;
or f0 (VV27V , d , c);
endmodule