module F1 (e , a , VV1V); 
input e , a;
output VV1V;
and f0 (VV1V , e , a);
endmodule