module F383 (VV381V , VV382V , VV383V); 
input VV381V , VV382V;
output VV383V;
and f0 (VV383V , VV381V , VV382V);
endmodule