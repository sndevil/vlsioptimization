module F113 (d , b , VV113V); 
input d , b;
output VV113V;
xor f0 (VV113V , d , b);
endmodule