module F173 (c , d , VV173V); 
input c , d;
output VV173V;
or f0 (VV173V , c , d);
endmodule