module F83 (e , d , VV83V); 
input e , d;
output VV83V;
xor f0 (VV83V , e , d);
endmodule