module F2 (VV1V , c , VV2V); 
input VV1V , c;
output VV2V;
and f0 (VV2V , VV1V , c);
endmodule