module F89 (c , d , VV89V); 
input c , d;
output VV89V;
and f0 (VV89V , c , d);
endmodule