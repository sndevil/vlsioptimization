module F240 (b , c , VV240V); 
input b , c;
output VV240V;
or f0 (VV240V , b , c);
endmodule