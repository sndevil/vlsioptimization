module F185 (VV183V , VV184V , VV185V); 
input VV183V , VV184V;
output VV185V;
or f0 (VV185V , VV183V , VV184V);
endmodule