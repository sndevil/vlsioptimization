module F353 (VV349V , VV352V , VV353V); 
input VV349V , VV352V;
output VV353V;
or f0 (VV353V , VV349V , VV352V);
endmodule