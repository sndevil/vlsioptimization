module F69 (a , b , VV69V); 
input a , b;
output VV69V;
xor f0 (VV69V , a , b);
endmodule