module F185 (e , a , VV185V); 
input e , a;
output VV185V;
or f0 (VV185V , e , a);
endmodule