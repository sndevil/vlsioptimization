module F2 (q , m , VV2V); 
input q , m;
output VV2V;
or f0 (VV2V , q , m);
endmodule