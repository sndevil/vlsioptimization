module F394 (VV362V , VV393V , VV394V); 
input VV362V , VV393V;
output VV394V;
or f0 (VV394V , VV362V , VV393V);
endmodule