module F343 (b , d , VV343V); 
input b , d;
output VV343V;
xor f0 (VV343V , b , d);
endmodule