module F73 (VV71V , VV72V , VV73V); 
input VV71V , VV72V;
output VV73V;
and f0 (VV73V , VV71V , VV72V);
endmodule