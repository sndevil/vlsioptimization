module F64 (VV62V , VV63V , VV64V); 
input VV62V , VV63V;
output VV64V;
xor f0 (VV64V , VV62V , VV63V);
endmodule