module F331 (VV299V , VV330V , VV331V); 
input VV299V , VV330V;
output VV331V;
or f0 (VV331V , VV299V , VV330V);
endmodule