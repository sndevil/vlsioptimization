module F138 (b , c , VV138V); 
input b , c;
output VV138V;
and f0 (VV138V , b , c);
endmodule