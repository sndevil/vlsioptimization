module F299 (VV283V , VV298V , VV299V); 
input VV283V , VV298V;
output VV299V;
or f0 (VV299V , VV283V , VV298V);
endmodule