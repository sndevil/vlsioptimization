module F39 (d , c , VV39V); 
input d , c;
output VV39V;
and f0 (VV39V , d , c);
endmodule