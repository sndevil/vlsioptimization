module F288 (a , b , VV288V); 
input a , b;
output VV288V;
or f0 (VV288V , a , b);
endmodule