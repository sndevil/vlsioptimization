module F161 (b , e , VV161V); 
input b , e;
output VV161V;
xor f0 (VV161V , b , e);
endmodule