module F187 (VV179V , VV186V , VV187V); 
input VV179V , VV186V;
output VV187V;
or f0 (VV187V , VV179V , VV186V);
endmodule