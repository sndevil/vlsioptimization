module F93 (VV89V , VV92V , VV93V); 
input VV89V , VV92V;
output VV93V;
or f0 (VV93V , VV89V , VV92V);
endmodule