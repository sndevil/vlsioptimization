module F19 (d , e , VV19V); 
input d , e;
output VV19V;
and f0 (VV19V , d , e);
endmodule