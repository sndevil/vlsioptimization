module F235 (VV219V , VV234V , VV235V); 
input VV219V , VV234V;
output VV235V;
and f0 (VV235V , VV219V , VV234V);
endmodule