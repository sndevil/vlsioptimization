module F294 (c , a , VV294V); 
input c , a;
output VV294V;
and f0 (VV294V , c , a);
endmodule