module F84 (VV82V , VV83V , VV84V); 
input VV82V , VV83V;
output VV84V;
xor f0 (VV84V , VV82V , VV83V);
endmodule