module F342 (e , b , VV342V); 
input e , b;
output VV342V;
xor f0 (VV342V , e , b);
endmodule