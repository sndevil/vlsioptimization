module F28 (VV26V , VV27V , VV28V); 
input VV26V , VV27V;
output VV28V;
xor f0 (VV28V , VV26V , VV27V);
endmodule