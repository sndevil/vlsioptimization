module F129 (d , a , VV129V); 
input d , a;
output VV129V;
xor f0 (VV129V , d , a);
endmodule