module F119 (VV117V , VV118V , VV119V); 
input VV117V , VV118V;
output VV119V;
or f0 (VV119V , VV117V , VV118V);
endmodule