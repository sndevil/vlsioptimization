module F119 (d , b , VV119V); 
input d , b;
output VV119V;
or f0 (VV119V , d , b);
endmodule