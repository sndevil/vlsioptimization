module F38 (d , a , VV38V); 
input d , a;
output VV38V;
wire WW37W0W;

not f0 (WW37W0W , d);
and f1 (VV38V , WW37W0W , a);
endmodule