module F310 (b , e , VV310V); 
input b , e;
output VV310V;
or f0 (VV310V , b , e);
endmodule