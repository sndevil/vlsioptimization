module F120 (VV118V , VV119V , VV120V); 
input VV118V , VV119V;
output VV120V;
xor f0 (VV120V , VV118V , VV119V);
endmodule