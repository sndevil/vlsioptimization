module F48 (b , d , VV48V); 
input b , d;
output VV48V;
xor f0 (VV48V , b , d);
endmodule