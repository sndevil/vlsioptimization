module F306 (VV302V , VV305V , VV306V); 
input VV302V , VV305V;
output VV306V;
and f0 (VV306V , VV302V , VV305V);
endmodule