module F91 (d , b , VV91V); 
input d , b;
output VV91V;
or f0 (VV91V , d , b);
endmodule