module F164 (b , a , VV164V); 
input b , a;
output VV164V;
and f0 (VV164V , b , a);
endmodule