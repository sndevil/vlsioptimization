module F123 (VV119V , VV122V , VV123V); 
input VV119V , VV122V;
output VV123V;
xor f0 (VV123V , VV119V , VV122V);
endmodule