module F260 (VV258V , VV259V , VV260V); 
input VV258V , VV259V;
output VV260V;
or f0 (VV260V , VV258V , VV259V);
endmodule