module F70 (b , e , VV70V); 
input b , e;
output VV70V;
and f0 (VV70V , b , e);
endmodule