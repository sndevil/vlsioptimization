module F43 (VV41V , VV42V , VV43V); 
input VV41V , VV42V;
output VV43V;
and f0 (VV43V , VV41V , VV42V);
endmodule