module F48 (d , a , VV48V); 
input d , a;
output VV48V;
or f0 (VV48V , d , a);
endmodule