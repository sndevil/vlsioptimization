module F45 (VV37V , VV44V , VV45V); 
input VV37V , VV44V;
output VV45V;
or f0 (VV45V , VV37V , VV44V);
endmodule