module F50 (d , a , VV50V); 
input d , a;
output VV50V;
xor f0 (VV50V , d , a);
endmodule