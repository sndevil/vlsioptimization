module F17 (b , c , VV17V); 
input b , c;
output VV17V;
xor f0 (VV17V , b , c);
endmodule