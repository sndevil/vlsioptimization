module F53 (VV49V , VV52V , VV53V); 
input VV49V , VV52V;
output VV53V;
or f0 (VV53V , VV49V , VV52V);
endmodule