module F45 (VV41V , VV44V , VV45V); 
input VV41V , VV44V;
output VV45V;
or f0 (VV45V , VV41V , VV44V);
endmodule