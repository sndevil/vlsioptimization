module F261 (b , d , VV261V); 
input b , d;
output VV261V;
and f0 (VV261V , b , d);
endmodule