module F208 (b , d , VV208V); 
input b , d;
output VV208V;
and f0 (VV208V , b , d);
endmodule