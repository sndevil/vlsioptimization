module F104 (VV102V , VV103V , VV104V); 
input VV102V , VV103V;
output VV104V;
or f0 (VV104V , VV102V , VV103V);
endmodule