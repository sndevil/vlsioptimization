module F183 (VV181V , VV182V , VV183V); 
input VV181V , VV182V;
output VV183V;
xor f0 (VV183V , VV181V , VV182V);
endmodule