module F38 (VV34V , VV37V , VV38V); 
input VV34V , VV37V;
output VV38V;
and f0 (VV38V , VV34V , VV37V);
endmodule