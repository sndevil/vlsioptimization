module F218 (VV214V , VV217V , VV218V); 
input VV214V , VV217V;
output VV218V;
and f0 (VV218V , VV214V , VV217V);
endmodule