module F220 (e , d , VV220V); 
input e , d;
output VV220V;
xor f0 (VV220V , e , d);
endmodule