module F386 (a , d , VV386V); 
input a , d;
output VV386V;
or f0 (VV386V , a , d);
endmodule