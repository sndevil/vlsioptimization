module F167 (a , c , VV167V); 
input a , c;
output VV167V;
xor f0 (VV167V , a , c);
endmodule