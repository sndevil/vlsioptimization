module F17 (b , e , VV17V); 
input b , e;
output VV17V;
and f0 (VV17V , b , e);
endmodule