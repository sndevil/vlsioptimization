module F23 (d , c , VV23V); 
input d , c;
output VV23V;
or f0 (VV23V , d , c);
endmodule