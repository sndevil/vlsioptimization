module F253 (VV251V , VV252V , VV253V); 
input VV251V , VV252V;
output VV253V;
xor f0 (VV253V , VV251V , VV252V);
endmodule