module F62 (b , d , VV62V); 
input b , d;
output VV62V;
or f0 (VV62V , b , d);
endmodule