module F108 (VV104V , VV107V , VV108V); 
input VV104V , VV107V;
output VV108V;
xor f0 (VV108V , VV104V , VV107V);
endmodule