module F88 (VV86V , VV87V , VV88V); 
input VV86V , VV87V;
output VV88V;
or f0 (VV88V , VV86V , VV87V);
endmodule