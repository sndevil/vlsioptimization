module F328 (VV324V , VV327V , VV328V); 
input VV324V , VV327V;
output VV328V;
and f0 (VV328V , VV324V , VV327V);
endmodule