module F117 (VV109V , VV116V , VV117V); 
input VV109V , VV116V;
output VV117V;
xor f0 (VV117V , VV109V , VV116V);
endmodule