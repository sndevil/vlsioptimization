module F15 (VV7V , VV14V , VV15V); 
input VV7V , VV14V;
output VV15V;
xor f0 (VV15V , VV7V , VV14V);
endmodule