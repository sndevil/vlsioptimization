module F369 (VV365V , VV368V , VV369V); 
input VV365V , VV368V;
output VV369V;
xor f0 (VV369V , VV365V , VV368V);
endmodule