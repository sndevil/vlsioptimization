module F37 (VV35V , VV36V , VV37V); 
input VV35V , VV36V;
output VV37V;
xor f0 (VV37V , VV35V , VV36V);
endmodule