module F114 (c , d , VV114V); 
input c , d;
output VV114V;
xor f0 (VV114V , c , d);
endmodule