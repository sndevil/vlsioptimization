module F149 (VV141V , VV148V , VV149V); 
input VV141V , VV148V;
output VV149V;
or f0 (VV149V , VV141V , VV148V);
endmodule