module F118 (c , b , VV118V); 
input c , b;
output VV118V;
xor f0 (VV118V , c , b);
endmodule