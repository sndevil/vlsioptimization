module F26 (b , d , VV26V); 
input b , d;
output VV26V;
xor f0 (VV26V , b , d);
endmodule