module F80 (b , a , VV80V); 
input b , a;
output VV80V;
and f0 (VV80V , b , a);
endmodule