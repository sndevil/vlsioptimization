module F116 (VV112V , VV115V , VV116V); 
input VV112V , VV115V;
output VV116V;
and f0 (VV116V , VV112V , VV115V);
endmodule