module F6 (a , c , VV6V); 
input a , c;
output VV6V;
xor f0 (VV6V , a , c);
endmodule