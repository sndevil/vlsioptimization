module F8 (b , d , VV8V); 
input b , d;
output VV8V;
or f0 (VV8V , b , d);
endmodule