module F62 (VV46V , VV61V , VV62V); 
input VV46V , VV61V;
output VV62V;
xor f0 (VV62V , VV46V , VV61V);
endmodule