module F135 (d , a , VV135V); 
input d , a;
output VV135V;
and f0 (VV135V , d , a);
endmodule