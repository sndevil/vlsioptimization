module F11 (e , b , VV11V); 
input e , b;
output VV11V;
or f0 (VV11V , e , b);
endmodule