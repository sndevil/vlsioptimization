module V1 (V#0#0# , a , c , V#1# , V#0#0# , q); 
