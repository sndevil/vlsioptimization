module F131 (b , c , VV131V); 
input b , c;
output VV131V;
or f0 (VV131V , b , c);
endmodule