module F380 (VV378V , VV379V , VV380V); 
input VV378V , VV379V;
output VV380V;
or f0 (VV380V , VV378V , VV379V);
endmodule