module F285 (e , a , VV285V); 
input e , a;
output VV285V;
or f0 (VV285V , e , a);
endmodule