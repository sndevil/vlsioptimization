module F86 (VV78V , VV85V , VV86V); 
input VV78V , VV85V;
output VV86V;
and f0 (VV86V , VV78V , VV85V);
endmodule