module F42 (b , d , VV42V); 
input b , d;
output VV42V;
or f0 (VV42V , b , d);
endmodule