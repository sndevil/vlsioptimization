module F360 (VV356V , VV359V , VV360V); 
input VV356V , VV359V;
output VV360V;
and f0 (VV360V , VV356V , VV359V);
endmodule