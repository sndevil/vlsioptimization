module F141 (VV127V , VV140V , VV141V); 
input VV127V , VV140V;
output VV141V;
or f0 (VV141V , VV127V , VV140V);
endmodule