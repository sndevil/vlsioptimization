module F8 (b , a , VV8V); 
input b , a;
output VV8V;
wire WW7W0W;

not f0 (WW7W0W , b);
and f1 (VV8V , a , WW7W0W);
endmodule