module F79 (e , d , VV79V); 
input e , d;
output VV79V;
or f0 (VV79V , e , d);
endmodule