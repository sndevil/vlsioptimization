module F176 (d , a , VV176V); 
input d , a;
output VV176V;
xor f0 (VV176V , d , a);
endmodule