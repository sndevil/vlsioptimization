module F151 (VV149V , VV150V , VV151V); 
input VV149V , VV150V;
output VV151V;
or f0 (VV151V , VV149V , VV150V);
endmodule