module F296 (VV294V , VV295V , VV296V); 
input VV294V , VV295V;
output VV296V;
or f0 (VV296V , VV294V , VV295V);
endmodule