module F87 (c , b , VV87V); 
input c , b;
output VV87V;
and f0 (VV87V , c , b);
endmodule