module F113 (e , a , VV113V); 
input e , a;
output VV113V;
and f0 (VV113V , e , a);
endmodule