module F18 (VV16V , VV17V , VV18V); 
input VV16V , VV17V;
output VV18V;
or f0 (VV18V , VV16V , VV17V);
endmodule