module F40 (e , b , VV40V); 
input e , b;
output VV40V;
xor f0 (VV40V , e , b);
endmodule