module F17 (d , c , VV17V); 
input d , c;
output VV17V;
and f0 (VV17V , d , c);
endmodule