module F211 (VV207V , VV210V , VV211V); 
input VV207V , VV210V;
output VV211V;
xor f0 (VV211V , VV207V , VV210V);
endmodule