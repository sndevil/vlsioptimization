module F180 (VV172V , VV179V , VV180V); 
input VV172V , VV179V;
output VV180V;
and f0 (VV180V , VV172V , VV179V);
endmodule