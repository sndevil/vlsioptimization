module F363 (a , b , VV363V); 
input a , b;
output VV363V;
or f0 (VV363V , a , b);
endmodule