module F234 (VV226V , VV233V , VV234V); 
input VV226V , VV233V;
output VV234V;
and f0 (VV234V , VV226V , VV233V);
endmodule