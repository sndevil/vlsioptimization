module F176 (d , b , VV176V); 
input d , b;
output VV176V;
or f0 (VV176V , d , b);
endmodule