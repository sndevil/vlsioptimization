module F221 (e , a , VV221V); 
input e , a;
output VV221V;
and f0 (VV221V , e , a);
endmodule