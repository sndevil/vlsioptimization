module F74 (VV72V , VV73V , VV74V); 
input VV72V , VV73V;
output VV74V;
and f0 (VV74V , VV72V , VV73V);
endmodule