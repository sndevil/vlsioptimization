module F19 (a , c , VV19V); 
input a , c;
output VV19V;
xor f0 (VV19V , a , c);
endmodule