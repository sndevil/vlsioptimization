module F132 (d , c , VV132V); 
input d , c;
output VV132V;
and f0 (VV132V , d , c);
endmodule