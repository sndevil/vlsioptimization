module F66 (VV64V , VV65V , VV66V); 
input VV64V , VV65V;
output VV66V;
and f0 (VV66V , VV64V , VV65V);
endmodule