module V2 (c , d , V#2#); 
input c , d;
output V#2#;
or f0 (V#2# , c , d);
endmodule