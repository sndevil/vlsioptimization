module F197 (VV165V , VV196V , VV197V); 
input VV165V , VV196V;
output VV197V;
or f0 (VV197V , VV165V , VV196V);
endmodule