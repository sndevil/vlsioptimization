module F141 (VV137V , VV140V , VV141V); 
input VV137V , VV140V;
output VV141V;
or f0 (VV141V , VV137V , VV140V);
endmodule