module F290 (VV286V , VV289V , VV290V); 
input VV286V , VV289V;
output VV290V;
or f0 (VV290V , VV286V , VV289V);
endmodule