module F373 (d , a , VV373V); 
input d , a;
output VV373V;
and f0 (VV373V , d , a);
endmodule