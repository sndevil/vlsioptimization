module F67 (e , b , VV67V); 
input e , b;
output VV67V;
or f0 (VV67V , e , b);
endmodule