module F352 (VV350V , VV351V , VV352V); 
input VV350V , VV351V;
output VV352V;
or f0 (VV352V , VV350V , VV351V);
endmodule