module F154 (d , e , VV154V); 
input d , e;
output VV154V;
and f0 (VV154V , d , e);
endmodule