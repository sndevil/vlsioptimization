module F304 (e , b , VV304V); 
input e , b;
output VV304V;
xor f0 (VV304V , e , b);
endmodule