module F74 (d , b , VV74V); 
input d , b;
output VV74V;
xor f0 (VV74V , d , b);
endmodule