module F73 (d , b , VV73V); 
input d , b;
output VV73V;
and f0 (VV73V , d , b);
endmodule