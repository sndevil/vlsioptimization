module F317 (VV315V , VV316V , VV317V); 
input VV315V , VV316V;
output VV317V;
and f0 (VV317V , VV315V , VV316V);
endmodule