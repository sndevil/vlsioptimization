module F148 (VV144V , VV147V , VV148V); 
input VV144V , VV147V;
output VV148V;
or f0 (VV148V , VV144V , VV147V);
endmodule