module F42 (d , e , VV42V); 
input d , e;
output VV42V;
or f0 (VV42V , d , e);
endmodule