module F271 (VV269V , VV270V , VV271V); 
input VV269V , VV270V;
output VV271V;
xor f0 (VV271V , VV269V , VV270V);
endmodule