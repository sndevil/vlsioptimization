module F94 (VV78V , VV93V , VV94V); 
input VV78V , VV93V;
output VV94V;
xor f0 (VV94V , VV78V , VV93V);
endmodule