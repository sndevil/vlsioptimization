module F181 (d , c , VV181V); 
input d , c;
output VV181V;
or f0 (VV181V , d , c);
endmodule