module F31 (e , b , VV31V); 
input e , b;
output VV31V;
or f0 (VV31V , e , b);
endmodule