module F158 (e , b , VV158V); 
input e , b;
output VV158V;
and f0 (VV158V , e , b);
endmodule