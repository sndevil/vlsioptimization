module F275 (VV271V , VV274V , VV275V); 
input VV271V , VV274V;
output VV275V;
or f0 (VV275V , VV271V , VV274V);
endmodule