module F55 (c , e , VV55V); 
input c , e;
output VV55V;
xor f0 (VV55V , c , e);
endmodule