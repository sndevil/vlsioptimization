module F242 (VV238V , VV241V , VV242V); 
input VV238V , VV241V;
output VV242V;
and f0 (VV242V , VV238V , VV241V);
endmodule