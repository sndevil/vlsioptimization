module F44 (VV40V , VV43V , VV44V); 
input VV40V , VV43V;
output VV44V;
and f0 (VV44V , VV40V , VV43V);
endmodule