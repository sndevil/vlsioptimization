module F111 (c , d , VV111V); 
input c , d;
output VV111V;
or f0 (VV111V , c , d);
endmodule