module F5 (q , i , VV5V); 
input q , i;
output VV5V;
and f0 (VV5V , q , i);
endmodule