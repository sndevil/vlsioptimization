module F382 (e , b , VV382V); 
input e , b;
output VV382V;
xor f0 (VV382V , e , b);
endmodule