module F86 (d , c , VV86V); 
input d , c;
output VV86V;
or f0 (VV86V , d , c);
endmodule