module F75 (VV71V , VV74V , VV75V); 
input VV71V , VV74V;
output VV75V;
xor f0 (VV75V , VV71V , VV74V);
endmodule