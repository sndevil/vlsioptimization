module F248 (VV246V , VV247V , VV248V); 
input VV246V , VV247V;
output VV248V;
or f0 (VV248V , VV246V , VV247V);
endmodule