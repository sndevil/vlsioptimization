module F41 (VV39V , VV40V , VV41V); 
input VV39V , VV40V;
output VV41V;
xor f0 (VV41V , VV39V , VV40V);
endmodule