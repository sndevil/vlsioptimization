module F170 (c , e , VV170V); 
input c , e;
output VV170V;
or f0 (VV170V , c , e);
endmodule