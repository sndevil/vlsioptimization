module F46 (VV38V , VV45V , VV46V); 
input VV38V , VV45V;
output VV46V;
and f0 (VV46V , VV38V , VV45V);
endmodule