module F90 (a , b , VV90V); 
input a , b;
output VV90V;
and f0 (VV90V , a , b);
endmodule