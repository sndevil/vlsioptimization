module F109 (VV105V , VV108V , VV109V); 
input VV105V , VV108V;
output VV109V;
or f0 (VV109V , VV105V , VV108V);
endmodule