module F153 (c , e , VV153V); 
input c , e;
output VV153V;
xor f0 (VV153V , c , e);
endmodule