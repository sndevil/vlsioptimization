module F103 (e , b , VV103V); 
input e , b;
output VV103V;
or f0 (VV103V , e , b);
endmodule