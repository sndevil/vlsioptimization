module F97 (a , b , VV97V); 
input a , b;
output VV97V;
and f0 (VV97V , a , b);
endmodule