module F157 (b , a , VV157V); 
input b , a;
output VV157V;
and f0 (VV157V , b , a);
endmodule