module F122 (a , d , VV122V); 
input a , d;
output VV122V;
xor f0 (VV122V , a , d);
endmodule