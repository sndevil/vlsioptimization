module F293 (VV291V , VV292V , VV293V); 
input VV291V , VV292V;
output VV293V;
or f0 (VV293V , VV291V , VV292V);
endmodule