module F341 (VV339V , VV340V , VV341V); 
input VV339V , VV340V;
output VV341V;
and f0 (VV341V , VV339V , VV340V);
endmodule