module F31 (b , a , VV31V); 
input b , a;
output VV31V;
xor f0 (VV31V , b , a);
endmodule