module F108 (VV106V , VV107V , VV108V); 
input VV106V , VV107V;
output VV108V;
and f0 (VV108V , VV106V , VV107V);
endmodule