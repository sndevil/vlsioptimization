module F297 (VV293V , VV296V , VV297V); 
input VV293V , VV296V;
output VV297V;
and f0 (VV297V , VV293V , VV296V);
endmodule