module F26 (e , d , VV26V); 
input e , d;
output VV26V;
or f0 (VV26V , e , d);
endmodule