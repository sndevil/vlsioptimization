module F41 (d , a , VV41V); 
input d , a;
output VV41V;
wire WW40W0W;

not f0 (WW40W0W , d);
and f1 (VV41V , a , WW40W0W);
endmodule