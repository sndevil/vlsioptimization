module F8 (b , a , VV8V); 
input b , a;
output VV8V;
or f0 (VV8V , b , a);
endmodule