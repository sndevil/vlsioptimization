module F63 (VV31V , VV62V , VV63V); 
input VV31V , VV62V;
output VV63V;
or f0 (VV63V , VV31V , VV62V);
endmodule