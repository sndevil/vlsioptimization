module F320 (VV318V , VV319V , VV320V); 
input VV318V , VV319V;
output VV320V;
or f0 (VV320V , VV318V , VV319V);
endmodule