module F76 (d , b , VV76V); 
input d , b;
output VV76V;
xor f0 (VV76V , d , b);
endmodule