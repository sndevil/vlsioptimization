module F255 (b , e , VV255V); 
input b , e;
output VV255V;
or f0 (VV255V , b , e);
endmodule