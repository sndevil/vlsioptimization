module F134 (VV102V , VV133V , VV134V); 
input VV102V , VV133V;
output VV134V;
and f0 (VV134V , VV102V , VV133V);
endmodule