module F334 (VV332V , VV333V , VV334V); 
input VV332V , VV333V;
output VV334V;
xor f0 (VV334V , VV332V , VV333V);
endmodule