module F69 (VV67V , VV68V , VV69V); 
input VV67V , VV68V;
output VV69V;
or f0 (VV69V , VV67V , VV68V);
endmodule