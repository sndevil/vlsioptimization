module F179 (VV175V , VV178V , VV179V); 
input VV175V , VV178V;
output VV179V;
or f0 (VV179V , VV175V , VV178V);
endmodule