module F63 (d , b , VV63V); 
input d , b;
output VV63V;
wire WW62W0W;

not f0 (WW62W0W , d);
or f1 (VV63V , WW62W0W , b);
endmodule