module F378 (c , d , VV378V); 
input c , d;
output VV378V;
and f0 (VV378V , c , d);
endmodule