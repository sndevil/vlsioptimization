module F47 (c , d , VV47V); 
input c , d;
output VV47V;
or f0 (VV47V , c , d);
endmodule