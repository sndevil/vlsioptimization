module F284 (a , b , VV284V); 
input a , b;
output VV284V;
or f0 (VV284V , a , b);
endmodule