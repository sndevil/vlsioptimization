module F32 (c , e , VV32V); 
input c , e;
output VV32V;
and f0 (VV32V , c , e);
endmodule