module F362 (VV346V , VV361V , VV362V); 
input VV346V , VV361V;
output VV362V;
or f0 (VV362V , VV346V , VV361V);
endmodule