module F228 (e , b , VV228V); 
input e , b;
output VV228V;
xor f0 (VV228V , e , b);
endmodule