module F78 (VV74V , VV77V , VV78V); 
input VV74V , VV77V;
output VV78V;
or f0 (VV78V , VV74V , VV77V);
endmodule