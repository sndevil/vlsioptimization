module F134 (VV130V , VV133V , VV134V); 
input VV130V , VV133V;
output VV134V;
or f0 (VV134V , VV130V , VV133V);
endmodule