module F156 (VV148V , VV155V , VV156V); 
input VV148V , VV155V;
output VV156V;
or f0 (VV156V , VV148V , VV155V);
endmodule