module F83 (d , a , VV83V); 
input d , a;
output VV83V;
or f0 (VV83V , d , a);
endmodule