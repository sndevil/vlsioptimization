module F292 (b , d , VV292V); 
input b , d;
output VV292V;
and f0 (VV292V , b , d);
endmodule