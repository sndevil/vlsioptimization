module F121 (e , c , VV121V); 
input e , c;
output VV121V;
or f0 (VV121V , e , c);
endmodule