module F93 (VV85V , VV92V , VV93V); 
input VV85V , VV92V;
output VV93V;
and f0 (VV93V , VV85V , VV92V);
endmodule