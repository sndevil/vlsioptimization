module F95 (b , e , VV95V); 
input b , e;
output VV95V;
and f0 (VV95V , b , e);
endmodule