module F111 (c , a , VV111V); 
input c , a;
output VV111V;
or f0 (VV111V , c , a);
endmodule