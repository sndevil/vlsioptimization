module F311 (c , d , VV311V); 
input c , d;
output VV311V;
xor f0 (VV311V , c , d);
endmodule