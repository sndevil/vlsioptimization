module F35 (c , b , VV35V); 
input c , b;
output VV35V;
or f0 (VV35V , c , b);
endmodule