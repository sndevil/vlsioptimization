module F183 (a , c , VV183V); 
input a , c;
output VV183V;
xor f0 (VV183V , a , c);
endmodule