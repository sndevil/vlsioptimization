module F146 (e , c , VV146V); 
input e , c;
output VV146V;
or f0 (VV146V , e , c);
endmodule