module F118 (d , c , VV118V); 
input d , c;
output VV118V;
or f0 (VV118V , d , c);
endmodule