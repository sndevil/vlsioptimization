module F128 (e , a , VV128V); 
input e , a;
output VV128V;
or f0 (VV128V , e , a);
endmodule