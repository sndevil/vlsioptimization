module F339 (e , b , VV339V); 
input e , b;
output VV339V;
xor f0 (VV339V , e , b);
endmodule