module F21 (VV19V , VV20V , VV21V); 
input VV19V , VV20V;
output VV21V;
xor f0 (VV21V , VV19V , VV20V);
endmodule