module F34 (b , d , VV34V); 
input b , d;
output VV34V;
or f0 (VV34V , b , d);
endmodule