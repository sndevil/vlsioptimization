module F4 (t , a , c , VV4V); 
input t , a , c;
output VV4V;
wire WW3W0W;

or f0 (WW3W0W , t , a);
and f1 (VV4V , WW3W0W , c);
endmodule