module F283 (VV275V , VV282V , VV283V); 
input VV275V , VV282V;
output VV283V;
and f0 (VV283V , VV275V , VV282V);
endmodule