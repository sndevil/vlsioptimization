module F188 (b , e , VV188V); 
input b , e;
output VV188V;
and f0 (VV188V , b , e);
endmodule