module F110 (a , b , VV110V); 
input a , b;
output VV110V;
and f0 (VV110V , a , b);
endmodule