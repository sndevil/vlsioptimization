module F350 (d , b , VV350V); 
input d , b;
output VV350V;
or f0 (VV350V , d , b);
endmodule