module F354 (d , e , VV354V); 
input d , e;
output VV354V;
xor f0 (VV354V , d , e);
endmodule