module F159 (VV157V , VV158V , VV159V); 
input VV157V , VV158V;
output VV159V;
and f0 (VV159V , VV157V , VV158V);
endmodule