module F54 (e , c , VV54V); 
input e , c;
output VV54V;
xor f0 (VV54V , e , c);
endmodule