module F236 (e , d , VV236V); 
input e , d;
output VV236V;
and f0 (VV236V , e , d);
endmodule