module F323 (c , d , VV323V); 
input c , d;
output VV323V;
xor f0 (VV323V , c , d);
endmodule