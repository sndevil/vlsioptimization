module F12 (d , a , VV12V); 
input d , a;
output VV12V;
or f0 (VV12V , d , a);
endmodule