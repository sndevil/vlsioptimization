module F39 (e , d , VV39V); 
input e , d;
output VV39V;
xor f0 (VV39V , e , d);
endmodule