module F1 (a , b , VV1V); 
input a , b;
output VV1V;
or f0 (VV1V , a , b);
endmodule