module F174 (a , c , VV174V); 
input a , c;
output VV174V;
or f0 (VV174V , a , c);
endmodule