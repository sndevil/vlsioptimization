module V2 (V#0#0# , a , b , V#1# , V#0#0# , c , a , V#1#0# , V#2# , V#1# , V#1#0#) 
