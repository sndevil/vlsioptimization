module F90 (e , a , VV90V); 
input e , a;
output VV90V;
and f0 (VV90V , e , a);
endmodule