module F286 (VV284V , VV285V , VV286V); 
input VV284V , VV285V;
output VV286V;
or f0 (VV286V , VV284V , VV285V);
endmodule