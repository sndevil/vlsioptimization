module F130 (VV128V , VV129V , VV130V); 
input VV128V , VV129V;
output VV130V;
or f0 (VV130V , VV128V , VV129V);
endmodule