module F332 (e , d , VV332V); 
input e , d;
output VV332V;
xor f0 (VV332V , e , d);
endmodule