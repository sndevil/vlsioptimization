module F77 (VV61V , VV76V , VV77V); 
input VV61V , VV76V;
output VV77V;
or f0 (VV77V , VV61V , VV76V);
endmodule