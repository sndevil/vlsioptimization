module F155 (VV153V , VV154V , VV155V); 
input VV153V , VV154V;
output VV155V;
or f0 (VV155V , VV153V , VV154V);
endmodule