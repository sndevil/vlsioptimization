module F351 (d , b , VV351V); 
input d , b;
output VV351V;
and f0 (VV351V , d , b);
endmodule