module F19 (d , b , VV19V); 
input d , b;
output VV19V;
wire WW18W0W;

not f0 (WW18W0W , d);
and f1 (VV19V , WW18W0W , b);
endmodule