module F47 (b , a , VV47V); 
input b , a;
output VV47V;
xor f0 (VV47V , b , a);
endmodule