module F156 (VV152V , VV155V , VV156V); 
input VV152V , VV155V;
output VV156V;
or f0 (VV156V , VV152V , VV155V);
endmodule