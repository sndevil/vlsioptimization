module F174 (c , d , VV174V); 
input c , d;
output VV174V;
and f0 (VV174V , c , d);
endmodule