module F26 (e , b , VV26V); 
input e , b;
output VV26V;
or f0 (VV26V , e , b);
endmodule