module F131 (VV127V , VV130V , VV131V); 
input VV127V , VV130V;
output VV131V;
and f0 (VV131V , VV127V , VV130V);
endmodule