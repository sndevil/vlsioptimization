module F358 (e , a , VV358V); 
input e , a;
output VV358V;
or f0 (VV358V , e , a);
endmodule