module F126 (VV94V , VV125V , VV126V); 
input VV94V , VV125V;
output VV126V;
and f0 (VV126V , VV94V , VV125V);
endmodule