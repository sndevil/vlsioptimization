module F34 (d , b , VV34V); 
input d , b;
output VV34V;
or f0 (VV34V , d , b);
endmodule