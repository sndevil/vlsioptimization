module F152 (VV150V , VV151V , VV152V); 
input VV150V , VV151V;
output VV152V;
and f0 (VV152V , VV150V , VV151V);
endmodule