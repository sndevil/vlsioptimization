module F245 (VV243V , VV244V , VV245V); 
input VV243V , VV244V;
output VV245V;
and f0 (VV245V , VV243V , VV244V);
endmodule