module F184 (b , e , VV184V); 
input b , e;
output VV184V;
xor f0 (VV184V , b , e);
endmodule