module F198 (c , e , VV198V); 
input c , e;
output VV198V;
and f0 (VV198V , c , e);
endmodule