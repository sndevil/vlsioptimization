module F72 (a , d , VV72V); 
input a , d;
output VV72V;
and f0 (VV72V , a , d);
endmodule