module F349 (VV347V , VV348V , VV349V); 
input VV347V , VV348V;
output VV349V;
or f0 (VV349V , VV347V , VV348V);
endmodule