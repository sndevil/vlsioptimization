module F177 (c , b , VV177V); 
input c , b;
output VV177V;
xor f0 (VV177V , c , b);
endmodule