module F168 (d , e , VV168V); 
input d , e;
output VV168V;
and f0 (VV168V , d , e);
endmodule