module F76 (VV68V , VV75V , VV76V); 
input VV68V , VV75V;
output VV76V;
xor f0 (VV76V , VV68V , VV75V);
endmodule