module F327 (VV325V , VV326V , VV327V); 
input VV325V , VV326V;
output VV327V;
or f0 (VV327V , VV325V , VV326V);
endmodule