module F345 (VV341V , VV344V , VV345V); 
input VV341V , VV344V;
output VV345V;
or f0 (VV345V , VV341V , VV344V);
endmodule