module F264 (VV260V , VV263V , VV264V); 
input VV260V , VV263V;
output VV264V;
or f0 (VV264V , VV260V , VV263V);
endmodule