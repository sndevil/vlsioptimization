module F344 (VV342V , VV343V , VV344V); 
input VV342V , VV343V;
output VV344V;
or f0 (VV344V , VV342V , VV343V);
endmodule