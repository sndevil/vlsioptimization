module F32 (b , d , VV32V); 
input b , d;
output VV32V;
or f0 (VV32V , b , d);
endmodule