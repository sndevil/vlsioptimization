module F142 (d , b , VV142V); 
input d , b;
output VV142V;
or f0 (VV142V , d , b);
endmodule