module F313 (VV309V , VV312V , VV313V); 
input VV309V , VV312V;
output VV313V;
or f0 (VV313V , VV309V , VV312V);
endmodule