module F181 (b , a , VV181V); 
input b , a;
output VV181V;
and f0 (VV181V , b , a);
endmodule