module F165 (VV149V , VV164V , VV165V); 
input VV149V , VV164V;
output VV165V;
and f0 (VV165V , VV149V , VV164V);
endmodule