module F95 (e , a , VV95V); 
input e , a;
output VV95V;
or f0 (VV95V , e , a);
endmodule