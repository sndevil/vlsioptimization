module F381 (d , c , VV381V); 
input d , c;
output VV381V;
or f0 (VV381V , d , c);
endmodule