module F125 (a , b , VV125V); 
input a , b;
output VV125V;
or f0 (VV125V , a , b);
endmodule