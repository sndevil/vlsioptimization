module F36 (c , a , VV36V); 
input c , a;
output VV36V;
and f0 (VV36V , c , a);
endmodule