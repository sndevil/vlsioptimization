module F178 (VV176V , VV177V , VV178V); 
input VV176V , VV177V;
output VV178V;
xor f0 (VV178V , VV176V , VV177V);
endmodule