module F50 (a , b , VV50V); 
input a , b;
output VV50V;
xor f0 (VV50V , a , b);
endmodule