module F182 (b , e , VV182V); 
input b , e;
output VV182V;
or f0 (VV182V , b , e);
endmodule