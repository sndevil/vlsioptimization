module F196 (VV180V , VV195V , VV196V); 
input VV180V , VV195V;
output VV196V;
and f0 (VV196V , VV180V , VV195V);
endmodule