module F295 (e , d , VV295V); 
input e , d;
output VV295V;
xor f0 (VV295V , e , d);
endmodule