module F145 (c , d , VV145V); 
input c , d;
output VV145V;
and f0 (VV145V , c , d);
endmodule