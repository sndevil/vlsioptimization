module F197 (VV195V , VV196V , VV197V); 
input VV195V , VV196V;
output VV197V;
xor f0 (VV197V , VV195V , VV196V);
endmodule