module F94 (e , c , VV94V); 
input e , c;
output VV94V;
and f0 (VV94V , e , c);
endmodule