module F209 (a , b , VV209V); 
input a , b;
output VV209V;
or f0 (VV209V , a , b);
endmodule