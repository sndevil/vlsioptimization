module F184 (a , b , VV184V); 
input a , b;
output VV184V;
xor f0 (VV184V , a , b);
endmodule