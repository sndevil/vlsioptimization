module F272 (b , a , VV272V); 
input b , a;
output VV272V;
xor f0 (VV272V , b , a);
endmodule