module F66 (a , c , VV66V); 
input a , c;
output VV66V;
xor f0 (VV66V , a , c);
endmodule