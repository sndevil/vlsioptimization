module F348 (e , b , VV348V); 
input e , b;
output VV348V;
or f0 (VV348V , e , b);
endmodule