module F251 (e , d , VV251V); 
input e , d;
output VV251V;
or f0 (VV251V , e , d);
endmodule