module F239 (c , d , VV239V); 
input c , d;
output VV239V;
or f0 (VV239V , c , d);
endmodule