module F196 (d , a , VV196V); 
input d , a;
output VV196V;
xor f0 (VV196V , d , a);
endmodule