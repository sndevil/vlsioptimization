module F189 (d , b , VV189V); 
input d , b;
output VV189V;
xor f0 (VV189V , d , b);
endmodule