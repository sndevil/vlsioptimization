module F3 (a , c , VV3V); 
input a , c;
output VV3V;
xor f0 (VV3V , a , c);
endmodule