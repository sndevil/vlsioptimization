module F241 (VV239V , VV240V , VV241V); 
input VV239V , VV240V;
output VV241V;
and f0 (VV241V , VV239V , VV240V);
endmodule