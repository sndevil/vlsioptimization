module F64 (e , c , VV64V); 
input e , c;
output VV64V;
or f0 (VV64V , e , c);
endmodule