module F146 (b , a , VV146V); 
input b , a;
output VV146V;
or f0 (VV146V , b , a);
endmodule