module F190 (VV188V , VV189V , VV190V); 
input VV188V , VV189V;
output VV190V;
xor f0 (VV190V , VV188V , VV189V);
endmodule