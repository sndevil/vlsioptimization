module F321 (VV317V , VV320V , VV321V); 
input VV317V , VV320V;
output VV321V;
or f0 (VV321V , VV317V , VV320V);
endmodule