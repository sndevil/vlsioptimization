module F51 (a , b , VV51V); 
input a , b;
output VV51V;
or f0 (VV51V , a , b);
endmodule