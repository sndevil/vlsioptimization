module F336 (e , d , VV336V); 
input e , d;
output VV336V;
or f0 (VV336V , e , d);
endmodule