module F203 (VV187V , VV202V , VV203V); 
input VV187V , VV202V;
output VV203V;
or f0 (VV203V , VV187V , VV202V);
endmodule