module F226 (VV222V , VV225V , VV226V); 
input VV222V , VV225V;
output VV226V;
and f0 (VV226V , VV222V , VV225V);
endmodule