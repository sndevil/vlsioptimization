module F92 (VV88V , VV91V , VV92V); 
input VV88V , VV91V;
output VV92V;
xor f0 (VV92V , VV88V , VV91V);
endmodule