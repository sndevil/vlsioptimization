module F165 (c , a , VV165V); 
input c , a;
output VV165V;
and f0 (VV165V , c , a);
endmodule