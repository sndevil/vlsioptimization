module F305 (VV303V , VV304V , VV305V); 
input VV303V , VV304V;
output VV305V;
or f0 (VV305V , VV303V , VV304V);
endmodule