module F36 (c , e , VV36V); 
input c , e;
output VV36V;
and f0 (VV36V , c , e);
endmodule