module F78 (VV46V , VV77V , VV78V); 
input VV46V , VV77V;
output VV78V;
and f0 (VV78V , VV46V , VV77V);
endmodule