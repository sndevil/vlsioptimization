module F325 (c , a , VV325V); 
input c , a;
output VV325V;
and f0 (VV325V , c , a);
endmodule