module F98 (a , c , VV98V); 
input a , c;
output VV98V;
or f0 (VV98V , a , c);
endmodule