module F63 (d , e , VV63V); 
input d , e;
output VV63V;
and f0 (VV63V , d , e);
endmodule