module F2 (a , b , VV2V); 
input a , b;
output VV2V;
or f0 (VV2V , a , b);
endmodule