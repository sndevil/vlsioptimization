module F281 (VV279V , VV280V , VV281V); 
input VV279V , VV280V;
output VV281V;
and f0 (VV281V , VV279V , VV280V);
endmodule