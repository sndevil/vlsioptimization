module F98 (d , a , VV98V); 
input d , a;
output VV98V;
xor f0 (VV98V , d , a);
endmodule