module F143 (a , d , VV143V); 
input a , d;
output VV143V;
xor f0 (VV143V , a , d);
endmodule