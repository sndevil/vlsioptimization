module F396 (VV268V' , VV395V , VV396V); 
input VV268V' , VV395V;
output VV396V;
and f0 (VV396V , VV268V' , VV395V);
endmodule