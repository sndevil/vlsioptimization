module F65 (e , d , VV65V); 
input e , d;
output VV65V;
xor f0 (VV65V , e , d);
endmodule