module F39 (d , a , VV39V); 
input d , a;
output VV39V;
and f0 (VV39V , d , a);
endmodule