module F125 (VV109V , VV124V , VV125V); 
input VV109V , VV124V;
output VV125V;
or f0 (VV125V , VV109V , VV124V);
endmodule