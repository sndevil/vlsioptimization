module F302 (VV300V , VV301V , VV302V); 
input VV300V , VV301V;
output VV302V;
or f0 (VV302V , VV300V , VV301V);
endmodule