module F379 (e , a , VV379V); 
input e , a;
output VV379V;
xor f0 (VV379V , e , a);
endmodule