module F206 (e , b , VV206V); 
input e , b;
output VV206V;
or f0 (VV206V , e , b);
endmodule