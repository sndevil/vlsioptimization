module F122 (VV120V , VV121V , VV122V); 
input VV120V , VV121V;
output VV122V;
and f0 (VV122V , VV120V , VV121V);
endmodule