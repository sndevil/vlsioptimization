module F73 (d , c , VV73V); 
input d , c;
output VV73V;
wire WW72W0W;

not f0 (WW72W0W , d);
and f1 (VV73V , WW72W0W , c);
endmodule