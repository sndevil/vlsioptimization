module F192 (c , b , VV192V); 
input c , b;
output VV192V;
or f0 (VV192V , c , b);
endmodule