module F329 (VV321V , VV328V , VV329V); 
input VV321V , VV328V;
output VV329V;
and f0 (VV329V , VV321V , VV328V);
endmodule