module F145 (c , b , VV145V); 
input c , b;
output VV145V;
or f0 (VV145V , c , b);
endmodule