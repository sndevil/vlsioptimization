module F133 (VV131V , VV132V , VV133V); 
input VV131V , VV132V;
output VV133V;
xor f0 (VV133V , VV131V , VV132V);
endmodule