module F96 (VV94V , VV95V , VV96V); 
input VV94V , VV95V;
output VV96V;
xor f0 (VV96V , VV94V , VV95V);
endmodule