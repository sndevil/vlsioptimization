module F300 (b , c , VV300V); 
input b , c;
output VV300V;
and f0 (VV300V , b , c);
endmodule