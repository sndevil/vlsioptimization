module F91 (VV89V , VV90V , VV91V); 
input VV89V , VV90V;
output VV91V;
xor f0 (VV91V , VV89V , VV90V);
endmodule