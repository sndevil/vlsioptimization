module F60 (VV56V , VV59V , VV60V); 
input VV56V , VV59V;
output VV60V;
xor f0 (VV60V , VV56V , VV59V);
endmodule