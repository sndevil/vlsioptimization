module F136 (b , a , VV136V); 
input b , a;
output VV136V;
xor f0 (VV136V , b , a);
endmodule