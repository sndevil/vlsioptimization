module F87 (c , b , VV87V); 
input c , b;
output VV87V;
xor f0 (VV87V , c , b);
endmodule