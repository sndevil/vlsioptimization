module F72 (d , e , VV72V); 
input d , e;
output VV72V;
or f0 (VV72V , d , e);
endmodule