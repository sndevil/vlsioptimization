module F9 (b , c , VV9V); 
input b , c;
output VV9V;
and f0 (VV9V , b , c);
endmodule