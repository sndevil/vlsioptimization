module F270 (d , c , VV270V); 
input d , c;
output VV270V;
xor f0 (VV270V , d , c);
endmodule