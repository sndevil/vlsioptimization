module F229 (VV227V , VV228V , VV229V); 
input VV227V , VV228V;
output VV229V;
and f0 (VV229V , VV227V , VV228V);
endmodule