module F324 (VV322V , VV323V , VV324V); 
input VV322V , VV323V;
output VV324V;
xor f0 (VV324V , VV322V , VV323V);
endmodule