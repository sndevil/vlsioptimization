module F26 (c , a , VV26V); 
input c , a;
output VV26V;
and f0 (VV26V , c , a);
endmodule