module F198 (VV134V , VV197V , VV198V); 
input VV134V , VV197V;
output VV198V;
xor f0 (VV198V , VV134V , VV197V);
endmodule