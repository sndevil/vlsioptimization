module F42 (a , b , VV42V); 
input a , b;
output VV42V;
xor f0 (VV42V , a , b);
endmodule