module F169 (VV167V , VV168V , VV169V); 
input VV167V , VV168V;
output VV169V;
or f0 (VV169V , VV167V , VV168V);
endmodule