module F166 (a , c , VV166V); 
input a , c;
output VV166V;
xor f0 (VV166V , a , c);
endmodule