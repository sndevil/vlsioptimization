module F58 (d , c , VV58V); 
input d , c;
output VV58V;
or f0 (VV58V , d , c);
endmodule