module F169 (a , e , VV169V); 
input a , e;
output VV169V;
or f0 (VV169V , a , e);
endmodule