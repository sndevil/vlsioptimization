module F51 (a , d , VV51V); 
input a , d;
output VV51V;
wire WW50W0W;

not f0 (WW50W0W , a);
or f1 (VV51V , WW50W0W , d);
endmodule