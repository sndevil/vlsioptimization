module F322 (c , d , VV322V); 
input c , d;
output VV322V;
and f0 (VV322V , c , d);
endmodule