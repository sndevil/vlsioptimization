module F27 (d , e , VV27V); 
input d , e;
output VV27V;
or f0 (VV27V , d , e);
endmodule