module F35 (c , d , VV35V); 
input c , d;
output VV35V;
xor f0 (VV35V , c , d);
endmodule