module F102 (a , d , VV102V); 
input a , d;
output VV102V;
or f0 (VV102V , a , d);
endmodule