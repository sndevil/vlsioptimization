module F57 (d , b , VV57V); 
input d , b;
output VV57V;
wire WW56W0W;

not f0 (WW56W0W , d);
and f1 (VV57V , b , WW56W0W);
endmodule