module F219 (VV211V , VV218V , VV219V); 
input VV211V , VV218V;
output VV219V;
and f0 (VV219V , VV211V , VV218V);
endmodule