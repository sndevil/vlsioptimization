module F35 (e , b , VV35V); 
input e , b;
output VV35V;
or f0 (VV35V , e , b);
endmodule