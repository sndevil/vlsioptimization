module F107 (d , c , VV107V); 
input d , c;
output VV107V;
or f0 (VV107V , d , c);
endmodule