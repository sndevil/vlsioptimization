module F252 (e , b , VV252V); 
input e , b;
output VV252V;
or f0 (VV252V , e , b);
endmodule