module F171 (VV169V , VV170V , VV171V); 
input VV169V , VV170V;
output VV171V;
xor f0 (VV171V , VV169V , VV170V);
endmodule