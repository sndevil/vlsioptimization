module F195 (d , a , VV195V); 
input d , a;
output VV195V;
and f0 (VV195V , d , a);
endmodule