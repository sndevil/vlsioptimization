module F223 (b , c , VV223V); 
input b , c;
output VV223V;
and f0 (VV223V , b , c);
endmodule