module F11 (c , e , VV11V); 
input c , e;
output VV11V;
xor f0 (VV11V , c , e);
endmodule