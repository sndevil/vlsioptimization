module F237 (c , d , VV237V); 
input c , d;
output VV237V;
xor f0 (VV237V , c , d);
endmodule