module F152 (b , d , VV152V); 
input b , d;
output VV152V;
xor f0 (VV152V , b , d);
endmodule