module F20 (c , d , VV20V); 
input c , d;
output VV20V;
and f0 (VV20V , c , d);
endmodule