module F42 (a , e , VV42V); 
input a , e;
output VV42V;
and f0 (VV42V , a , e);
endmodule