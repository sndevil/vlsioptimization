module F1 (k , e , VV1V); 
input k , e;
output VV1V;
xor f0 (VV1V , k , e);
endmodule