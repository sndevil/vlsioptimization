module F333 (a , e , VV333V); 
input a , e;
output VV333V;
xor f0 (VV333V , a , e);
endmodule