module F85 (VV81V , VV84V , VV85V); 
input VV81V , VV84V;
output VV85V;
and f0 (VV85V , VV81V , VV84V);
endmodule