module F57 (e , b , VV57V); 
input e , b;
output VV57V;
xor f0 (VV57V , e , b);
endmodule