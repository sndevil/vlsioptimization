module F16 (c , d , VV16V); 
input c , d;
output VV16V;
and f0 (VV16V , c , d);
endmodule