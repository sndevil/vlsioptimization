module F126 (a , c , VV126V); 
input a , c;
output VV126V;
and f0 (VV126V , a , c);
endmodule