module F346 (VV338V , VV345V , VV346V); 
input VV338V , VV345V;
output VV346V;
xor f0 (VV346V , VV338V , VV345V);
endmodule