module F212 (c , b , VV212V); 
input c , b;
output VV212V;
and f0 (VV212V , c , b);
endmodule