module F289 (VV287V , VV288V , VV289V); 
input VV287V , VV288V;
output VV289V;
and f0 (VV289V , VV287V , VV288V);
endmodule