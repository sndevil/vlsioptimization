module F188 (b , d , VV188V); 
input b , d;
output VV188V;
and f0 (VV188V , b , d);
endmodule