module F17 (a , e , VV17V); 
input a , e;
output VV17V;
xor f0 (VV17V , a , e);
endmodule