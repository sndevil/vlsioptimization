module F33 (a , c , VV33V); 
input a , c;
output VV33V;
and f0 (VV33V , a , c);
endmodule