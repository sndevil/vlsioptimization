module F96 (e , a , VV96V); 
input e , a;
output VV96V;
or f0 (VV96V , e , a);
endmodule