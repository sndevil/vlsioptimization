module F (VV1V); 
;
output VV1V;
endmodule