module F41 (e , d , VV41V); 
input e , d;
output VV41V;
or f0 (VV41V , e , d);
endmodule