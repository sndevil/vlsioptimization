module F43 (e , c , VV43V); 
input e , c;
output VV43V;
and f0 (VV43V , e , c);
endmodule