module F175 (VV173V , VV174V , VV175V); 
input VV173V , VV174V;
output VV175V;
and f0 (VV175V , VV173V , VV174V);
endmodule