module F67 (c , d , VV67V); 
input c , d;
output VV67V;
and f0 (VV67V , c , d);
endmodule