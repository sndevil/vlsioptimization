module F157 (a , c , VV157V); 
input a , c;
output VV157V;
or f0 (VV157V , a , c);
endmodule