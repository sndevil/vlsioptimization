module F167 (d , a , VV167V); 
input d , a;
output VV167V;
xor f0 (VV167V , d , a);
endmodule