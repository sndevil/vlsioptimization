module F44 (VV42V , VV43V , VV44V); 
input VV42V , VV43V;
output VV44V;
or f0 (VV44V , VV42V , VV43V);
endmodule