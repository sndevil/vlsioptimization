module F357 (d , a , VV357V); 
input d , a;
output VV357V;
xor f0 (VV357V , d , a);
endmodule