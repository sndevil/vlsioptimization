module F4 (d , a , VV4V); 
input d , a;
output VV4V;
wire WW3W0W;

not f0 (WW3W0W , d);
and f1 (VV4V , a , WW3W0W);
endmodule