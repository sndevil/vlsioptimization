module F23 (b , c , VV23V); 
input b , c;
output VV23V;
and f0 (VV23V , b , c);
endmodule