module F192 (c , d , VV192V); 
input c , d;
output VV192V;
xor f0 (VV192V , c , d);
endmodule