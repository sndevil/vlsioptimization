module F194 (VV190V , VV193V , VV194V); 
input VV190V , VV193V;
output VV194V;
xor f0 (VV194V , VV190V , VV193V);
endmodule