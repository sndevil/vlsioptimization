module F375 (VV373V , VV374V , VV375V); 
input VV373V , VV374V;
output VV375V;
xor f0 (VV375V , VV373V , VV374V);
endmodule