module F199 (e , d , VV199V); 
input e , d;
output VV199V;
or f0 (VV199V , e , d);
endmodule