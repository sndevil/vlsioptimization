module F180 (b , c , VV180V); 
input b , c;
output VV180V;
and f0 (VV180V , b , c);
endmodule