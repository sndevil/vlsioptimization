module F168 (VV166V , VV167V , VV168V); 
input VV166V , VV167V;
output VV168V;
xor f0 (VV168V , VV166V , VV167V);
endmodule