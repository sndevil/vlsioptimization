module F389 (c , a , VV389V); 
input c , a;
output VV389V;
and f0 (VV389V , c , a);
endmodule