module F262 (b , e , VV262V); 
input b , e;
output VV262V;
or f0 (VV262V , b , e);
endmodule