module F200 (VV198V , VV199V , VV200V); 
input VV198V , VV199V;
output VV200V;
and f0 (VV200V , VV198V , VV199V);
endmodule