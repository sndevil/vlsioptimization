module F172 (VV168V , VV171V , VV172V); 
input VV168V , VV171V;
output VV172V;
or f0 (VV172V , VV168V , VV171V);
endmodule