module F268 (VV204V , VV267V , VV268V); 
input VV204V , VV267V;
output VV268V;
or f0 (VV268V , VV204V , VV267V);
endmodule