module F247 (b , c , VV247V); 
input b , c;
output VV247V;
or f0 (VV247V , b , c);
endmodule