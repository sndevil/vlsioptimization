module F191 (b , d , VV191V); 
input b , d;
output VV191V;
and f0 (VV191V , b , d);
endmodule