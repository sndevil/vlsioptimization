module F187 (VV183V , VV186V , VV187V); 
input VV183V , VV186V;
output VV187V;
or f0 (VV187V , VV183V , VV186V);
endmodule