module F4 (t , b , VV4V); 
input t , b;
output VV4V;
wire WW3W0W;

not f0 (WW3W0W , t);
or f1 (VV4V , b , WW3W0W);
endmodule