module F368 (VV366V , VV367V , VV368V); 
input VV366V , VV367V;
output VV368V;
and f0 (VV368V , VV366V , VV367V);
endmodule