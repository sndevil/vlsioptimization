module F58 (d , a , VV58V); 
input d , a;
output VV58V;
or f0 (VV58V , d , a);
endmodule