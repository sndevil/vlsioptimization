module F366 (b , e , VV366V); 
input b , e;
output VV366V;
xor f0 (VV366V , b , e);
endmodule