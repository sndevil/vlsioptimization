module F115 (VV113V , VV114V , VV115V); 
input VV113V , VV114V;
output VV115V;
and f0 (VV115V , VV113V , VV114V);
endmodule