module F265 (VV257V , VV264V , VV265V); 
input VV257V , VV264V;
output VV265V;
or f0 (VV265V , VV257V , VV264V);
endmodule