module F233 (VV229V , VV232V , VV233V); 
input VV229V , VV232V;
output VV233V;
and f0 (VV233V , VV229V , VV232V);
endmodule