module F355 (c , d , VV355V); 
input c , d;
output VV355V;
xor f0 (VV355V , c , d);
endmodule