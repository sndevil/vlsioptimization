module F338 (VV334V , VV337V , VV338V); 
input VV334V , VV337V;
output VV338V;
or f0 (VV338V , VV334V , VV337V);
endmodule