module F67 (VV65V , VV66V , VV67V); 
input VV65V , VV66V;
output VV67V;
xor f0 (VV67V , VV65V , VV66V);
endmodule