module F376 (VV372V , VV375V , VV376V); 
input VV372V , VV375V;
output VV376V;
and f0 (VV376V , VV372V , VV375V);
endmodule