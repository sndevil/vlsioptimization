module F326 (b , e , VV326V); 
input b , e;
output VV326V;
and f0 (VV326V , b , e);
endmodule