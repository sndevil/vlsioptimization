module F390 (VV388V , VV389V , VV390V); 
input VV388V , VV389V;
output VV390V;
and f0 (VV390V , VV388V , VV389V);
endmodule