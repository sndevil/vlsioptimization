module F371 (e , c , VV371V); 
input e , c;
output VV371V;
xor f0 (VV371V , e , c);
endmodule