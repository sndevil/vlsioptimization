module F356 (VV354V , VV355V , VV356V); 
input VV354V , VV355V;
output VV356V;
or f0 (VV356V , VV354V , VV355V);
endmodule