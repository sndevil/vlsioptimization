module F115 (VV113V , VV114V , VV115V); 
input VV113V , VV114V;
output VV115V;
xor f0 (VV115V , VV113V , VV114V);
endmodule