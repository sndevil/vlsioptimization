module F199 (VV71V , VV198V , VV199V); 
input VV71V , VV198V;
output VV199V;
xor f0 (VV199V , VV71V , VV198V);
endmodule