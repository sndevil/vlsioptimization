module F64 (a , b , VV64V); 
input a , b;
output VV64V;
and f0 (VV64V , a , b);
endmodule