module F72 (e , d , VV72V); 
input e , d;
output VV72V;
xor f0 (VV72V , e , d);
endmodule