module F24 (a , e , VV24V); 
input a , e;
output VV24V;
or f0 (VV24V , a , e);
endmodule