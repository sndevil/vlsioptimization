module F2 (j , h , VV2V); 
input j , h;
output VV2V;
and f0 (VV2V , j , h);
endmodule