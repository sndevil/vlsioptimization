module F301 (a , b , VV301V); 
input a , b;
output VV301V;
or f0 (VV301V , a , b);
endmodule