module F149 (e , d , VV149V); 
input e , d;
output VV149V;
or f0 (VV149V , e , d);
endmodule