module F11 (d , e , VV11V); 
input d , e;
output VV11V;
and f0 (VV11V , d , e);
endmodule