module F315 (a , d , VV315V); 
input a , d;
output VV315V;
xor f0 (VV315V , a , d);
endmodule