module F132 (VV124V , VV131V , VV132V); 
input VV124V , VV131V;
output VV132V;
and f0 (VV132V , VV124V , VV131V);
endmodule