module F372 (VV370V , VV371V , VV372V); 
input VV370V , VV371V;
output VV372V;
or f0 (VV372V , VV370V , VV371V);
endmodule