module F (VV2V); 
;
output VV2V;
endmodule