module V1 (b , a , V#1#); 
input b , a;
output V#1#;
wire W#0#0#;

not f0 (W#0#0# , b);
and f1 (V#1# , W#0#0# , a);
endmodule