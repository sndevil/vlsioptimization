module F377 (VV369V , VV376V , VV377V); 
input VV369V , VV376V;
output VV377V;
or f0 (VV377V , VV369V , VV376V);
endmodule