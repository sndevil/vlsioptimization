module F48 (e , c , VV48V); 
input e , c;
output VV48V;
and f0 (VV48V , e , c);
endmodule