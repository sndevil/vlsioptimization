module F65 (b , a , VV65V); 
input b , a;
output VV65V;
or f0 (VV65V , b , a);
endmodule