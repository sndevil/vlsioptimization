module F43 (e , b , VV43V); 
input e , b;
output VV43V;
and f0 (VV43V , e , b);
endmodule