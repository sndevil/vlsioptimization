module F57 (a , d , VV57V); 
input a , d;
output VV57V;
and f0 (VV57V , a , d);
endmodule