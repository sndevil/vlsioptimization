module F318 (b , c , VV318V); 
input b , c;
output VV318V;
and f0 (VV318V , b , c);
endmodule