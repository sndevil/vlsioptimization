module F123 (VV121V , VV122V , VV123V); 
input VV121V , VV122V;
output VV123V;
and f0 (VV123V , VV121V , VV122V);
endmodule