module F150 (b , e , VV150V); 
input b , e;
output VV150V;
xor f0 (VV150V , b , e);
endmodule