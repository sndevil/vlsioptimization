module F107 (VV105V , VV106V , VV107V); 
input VV105V , VV106V;
output VV107V;
xor f0 (VV107V , VV105V , VV106V);
endmodule