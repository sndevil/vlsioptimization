module F37 (VV33V , VV36V , VV37V); 
input VV33V , VV36V;
output VV37V;
and f0 (VV37V , VV33V , VV36V);
endmodule