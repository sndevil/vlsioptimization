module F71 (d , e , VV71V); 
input d , e;
output VV71V;
and f0 (VV71V , d , e);
endmodule