module F337 (VV335V , VV336V , VV337V); 
input VV335V , VV336V;
output VV337V;
xor f0 (VV337V , VV335V , VV336V);
endmodule