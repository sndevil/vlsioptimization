module F263 (VV261V , VV262V , VV263V); 
input VV261V , VV262V;
output VV263V;
xor f0 (VV263V , VV261V , VV262V);
endmodule