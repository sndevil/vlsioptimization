module F274 (VV272V , VV273V , VV274V); 
input VV272V , VV273V;
output VV274V;
and f0 (VV274V , VV272V , VV273V);
endmodule