module F12 (d , e , VV12V); 
input d , e;
output VV12V;
xor f0 (VV12V , d , e);
endmodule