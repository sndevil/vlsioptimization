module F55 (a , d , VV55V); 
input a , d;
output VV55V;
xor f0 (VV55V , a , d);
endmodule