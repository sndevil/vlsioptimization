module F249 (VV245V , VV248V , VV249V); 
input VV245V , VV248V;
output VV249V;
xor f0 (VV249V , VV245V , VV248V);
endmodule