module F82 (b , a , VV82V); 
input b , a;
output VV82V;
and f0 (VV82V , b , a);
endmodule