module F280 (b , e , VV280V); 
input b , e;
output VV280V;
and f0 (VV280V , b , e);
endmodule