module F47 (b , c , VV47V); 
input b , c;
output VV47V;
and f0 (VV47V , b , c);
endmodule