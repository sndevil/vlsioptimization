module F347 (d , a , VV347V); 
input d , a;
output VV347V;
and f0 (VV347V , d , a);
endmodule