module F231 (b , c , VV231V); 
input b , c;
output VV231V;
xor f0 (VV231V , b , c);
endmodule