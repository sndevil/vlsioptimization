module F279 (b , d , VV279V); 
input b , d;
output VV279V;
and f0 (VV279V , b , d);
endmodule