module F68 (e , a , VV68V); 
input e , a;
output VV68V;
and f0 (VV68V , e , a);
endmodule