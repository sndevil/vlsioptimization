module F170 (VV166V , VV169V , VV170V); 
input VV166V , VV169V;
output VV170V;
xor f0 (VV170V , VV166V , VV169V);
endmodule