module F101 (VV97V , VV100V , VV101V); 
input VV97V , VV100V;
output VV101V;
xor f0 (VV101V , VV97V , VV100V);
endmodule