module F137 (VV135V , VV136V , VV137V); 
input VV135V , VV136V;
output VV137V;
or f0 (VV137V , VV135V , VV136V);
endmodule