module F191 (c , d , VV191V); 
input c , d;
output VV191V;
or f0 (VV191V , c , d);
endmodule