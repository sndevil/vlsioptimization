module F8 (d , a , VV8V); 
input d , a;
output VV8V;
xor f0 (VV8V , d , a);
endmodule