module F307 (d , c , VV307V); 
input d , c;
output VV307V;
xor f0 (VV307V , d , c);
endmodule