module F27 (b , e , VV27V); 
input b , e;
output VV27V;
or f0 (VV27V , b , e);
endmodule