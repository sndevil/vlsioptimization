module F207 (VV205V , VV206V , VV207V); 
input VV205V , VV206V;
output VV207V;
or f0 (VV207V , VV205V , VV206V);
endmodule