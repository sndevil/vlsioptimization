module F88 (c , a , VV88V); 
input c , a;
output VV88V;
or f0 (VV88V , c , a);
endmodule