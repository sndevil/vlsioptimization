module F154 (VV152V , VV153V , VV154V); 
input VV152V , VV153V;
output VV154V;
and f0 (VV154V , VV152V , VV153V);
endmodule