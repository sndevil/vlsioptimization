module F161 (e , c , VV161V); 
input e , c;
output VV161V;
and f0 (VV161V , e , c);
endmodule