module F365 (VV363V , VV364V , VV365V); 
input VV363V , VV364V;
output VV365V;
and f0 (VV365V , VV363V , VV364V);
endmodule