module F144 (VV142V , VV143V , VV144V); 
input VV142V , VV143V;
output VV144V;
or f0 (VV144V , VV142V , VV143V);
endmodule