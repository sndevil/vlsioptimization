module F16 (d , a , VV16V); 
input d , a;
output VV16V;
or f0 (VV16V , d , a);
endmodule