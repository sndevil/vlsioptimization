module F75 (b , c , VV75V); 
input b , c;
output VV75V;
and f0 (VV75V , b , c);
endmodule