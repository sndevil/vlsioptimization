module F225 (VV223V , VV224V , VV225V); 
input VV223V , VV224V;
output VV225V;
or f0 (VV225V , VV223V , VV224V);
endmodule