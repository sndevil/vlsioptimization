module F81 (VV79V , VV80V , VV81V); 
input VV79V , VV80V;
output VV81V;
or f0 (VV81V , VV79V , VV80V);
endmodule