module F215 (d , b , VV215V); 
input d , b;
output VV215V;
or f0 (VV215V , d , b);
endmodule