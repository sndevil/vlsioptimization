module F278 (VV276V , VV277V , VV278V); 
input VV276V , VV277V;
output VV278V;
or f0 (VV278V , VV276V , VV277V);
endmodule