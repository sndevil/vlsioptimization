module F59 (VV57V , VV58V , VV59V); 
input VV57V , VV58V;
output VV59V;
or f0 (VV59V , VV57V , VV58V);
endmodule