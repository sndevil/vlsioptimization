module F140 (VV138V , VV139V , VV140V); 
input VV138V , VV139V;
output VV140V;
and f0 (VV140V , VV138V , VV139V);
endmodule