module F2 (b , e , VV2V); 
input b , e;
output VV2V;
xor f0 (VV2V , b , e);
endmodule