module F105 (e , d , VV105V); 
input e , d;
output VV105V;
xor f0 (VV105V , e , d);
endmodule