module F177 (e , b , VV177V); 
input e , b;
output VV177V;
and f0 (VV177V , e , b);
endmodule