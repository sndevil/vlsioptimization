module F153 (b , d , VV153V); 
input b , d;
output VV153V;
and f0 (VV153V , b , d);
endmodule