module F238 (VV236V , VV237V , VV238V); 
input VV236V , VV237V;
output VV238V;
or f0 (VV238V , VV236V , VV237V);
endmodule