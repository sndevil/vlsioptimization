module F173 (e , d , VV173V); 
input e , d;
output VV173V;
or f0 (VV173V , e , d);
endmodule