module F244 (c , e , VV244V); 
input c , e;
output VV244V;
or f0 (VV244V , c , e);
endmodule