module F56 (VV54V , VV55V , VV56V); 
input VV54V , VV55V;
output VV56V;
or f0 (VV56V , VV54V , VV55V);
endmodule