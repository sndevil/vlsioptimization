module F58 (c , a , VV58V); 
input c , a;
output VV58V;
wire WW57W0W;

not f0 (WW57W0W , c);
and f1 (VV58V , WW57W0W , a);
endmodule