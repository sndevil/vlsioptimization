module F9 (a , d , VV9V); 
input a , d;
output VV9V;
and f0 (VV9V , a , d);
endmodule