module F106 (c , a , VV106V); 
input c , a;
output VV106V;
or f0 (VV106V , c , a);
endmodule