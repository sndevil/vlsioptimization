module F20 (c , d , VV20V); 
input c , d;
output VV20V;
wire WW19W0W;

not f0 (WW19W0W , c);
and f1 (VV20V , WW19W0W , d);
endmodule