module F258 (a , b , VV258V); 
input a , b;
output VV258V;
and f0 (VV258V , a , b);
endmodule