module F163 (VV159V , VV162V , VV163V); 
input VV159V , VV162V;
output VV163V;
xor f0 (VV163V , VV159V , VV162V);
endmodule