module F312 (VV310V , VV311V , VV312V); 
input VV310V , VV311V;
output VV312V;
or f0 (VV312V , VV310V , VV311V);
endmodule