module F89 (VV87V , VV88V , VV89V); 
input VV87V , VV88V;
output VV89V;
and f0 (VV89V , VV87V , VV88V);
endmodule