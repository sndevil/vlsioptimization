module F164 (VV156V , VV163V , VV164V); 
input VV156V , VV163V;
output VV164V;
and f0 (VV164V , VV156V , VV163V);
endmodule