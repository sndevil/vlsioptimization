module F124 (VV116V , VV123V , VV124V); 
input VV116V , VV123V;
output VV124V;
and f0 (VV124V , VV116V , VV123V);
endmodule