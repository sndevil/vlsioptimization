module F186 (VV184V , VV185V , VV186V); 
input VV184V , VV185V;
output VV186V;
and f0 (VV186V , VV184V , VV185V);
endmodule