module F139 (VV137V , VV138V , VV139V); 
input VV137V , VV138V;
output VV139V;
and f0 (VV139V , VV137V , VV138V);
endmodule