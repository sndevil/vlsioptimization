module F385 (a , d , VV385V); 
input a , d;
output VV385V;
xor f0 (VV385V , a , d);
endmodule