module F139 (a , e , VV139V); 
input a , e;
output VV139V;
xor f0 (VV139V , a , e);
endmodule