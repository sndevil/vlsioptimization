module F133 (VV117V , VV132V , VV133V); 
input VV117V , VV132V;
output VV133V;
or f0 (VV133V , VV117V , VV132V);
endmodule