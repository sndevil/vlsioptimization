module F316 (d , e , VV316V); 
input d , e;
output VV316V;
and f0 (VV316V , d , e);
endmodule