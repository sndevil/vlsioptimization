module F309 (VV307V , VV308V , VV309V); 
input VV307V , VV308V;
output VV309V;
xor f0 (VV309V , VV307V , VV308V);
endmodule