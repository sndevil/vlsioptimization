module F40 (d , c , VV40V); 
input d , c;
output VV40V;
xor f0 (VV40V , d , c);
endmodule