module F24 (c , e , VV24V); 
input c , e;
output VV24V;
or f0 (VV24V , c , e);
endmodule