module F182 (VV180V , VV181V , VV182V); 
input VV180V , VV181V;
output VV182V;
or f0 (VV182V , VV180V , VV181V);
endmodule