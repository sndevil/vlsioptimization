module F254 (c , a , VV254V); 
input c , a;
output VV254V;
and f0 (VV254V , c , a);
endmodule