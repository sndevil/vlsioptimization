module F387 (VV385V , VV386V , VV387V); 
input VV385V , VV386V;
output VV387V;
or f0 (VV387V , VV385V , VV386V);
endmodule