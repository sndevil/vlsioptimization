module F58 (a , e , VV58V); 
input a , e;
output VV58V;
and f0 (VV58V , a , e);
endmodule