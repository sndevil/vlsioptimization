module F77 (VV73V , VV76V , VV77V); 
input VV73V , VV76V;
output VV77V;
and f0 (VV77V , VV73V , VV76V);
endmodule