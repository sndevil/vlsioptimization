module F155 (VV151V , VV154V , VV155V); 
input VV151V , VV154V;
output VV155V;
and f0 (VV155V , VV151V , VV154V);
endmodule