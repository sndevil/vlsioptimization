module F276 (d , a , VV276V); 
input d , a;
output VV276V;
xor f0 (VV276V , d , a);
endmodule