module F340 (d , e , VV340V); 
input d , e;
output VV340V;
xor f0 (VV340V , d , e);
endmodule