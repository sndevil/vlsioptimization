module F10 (VV8V , VV9V , VV10V); 
input VV8V , VV9V;
output VV10V;
or f0 (VV10V , VV8V , VV9V);
endmodule