module F38 (a , b , VV38V); 
input a , b;
output VV38V;
xor f0 (VV38V , a , b);
endmodule