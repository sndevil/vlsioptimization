module F202 (VV194V , VV201V , VV202V); 
input VV194V , VV201V;
output VV202V;
or f0 (VV202V , VV194V , VV201V);
endmodule