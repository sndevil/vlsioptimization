module F367 (d , c , VV367V); 
input d , c;
output VV367V;
and f0 (VV367V , d , c);
endmodule