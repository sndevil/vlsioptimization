module F213 (b , a , VV213V); 
input b , a;
output VV213V;
or f0 (VV213V , b , a);
endmodule