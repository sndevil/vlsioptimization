module F70 (VV66V , VV69V , VV70V); 
input VV66V , VV69V;
output VV70V;
or f0 (VV70V , VV66V , VV69V);
endmodule