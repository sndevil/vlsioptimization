module F4 (d , a , VV4V); 
input d , a;
output VV4V;
xor f0 (VV4V , d , a);
endmodule