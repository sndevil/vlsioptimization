module F319 (d , b , VV319V); 
input d , b;
output VV319V;
and f0 (VV319V , d , b);
endmodule