module F397 (VV141V , VV396V , VV397V); 
input VV141V , VV396V;
output VV397V;
xor f0 (VV397V , VV141V , VV396V);
endmodule