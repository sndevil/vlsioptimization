module F79 (c , a , VV79V); 
input c , a;
output VV79V;
and f0 (VV79V , c , a);
endmodule