module F205 (b , c , VV205V); 
input b , c;
output VV205V;
or f0 (VV205V , b , c);
endmodule