module F65 (d , c , VV65V); 
input d , c;
output VV65V;
or f0 (VV65V , d , c);
endmodule