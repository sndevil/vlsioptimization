module F224 (a , b , VV224V); 
input a , b;
output VV224V;
and f0 (VV224V , a , b);
endmodule