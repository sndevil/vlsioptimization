module F4 (c , m , VV4V); 
input c , m;
output VV4V;
or f0 (VV4V , c , m);
endmodule