module F193 (VV191V , VV192V , VV193V); 
input VV191V , VV192V;
output VV193V;
xor f0 (VV193V , VV191V , VV192V);
endmodule