module F82 (c , e , VV82V); 
input c , e;
output VV82V;
xor f0 (VV82V , c , e);
endmodule