module F140 (VV134V , VV139V , VV140V); 
input VV134V , VV139V;
output VV140V;
xor f0 (VV140V , VV134V , VV139V);
endmodule