module F7 (VV5V , VV6V , VV7V); 
input VV5V , VV6V;
output VV7V;
and f0 (VV7V , VV5V , VV6V);
endmodule