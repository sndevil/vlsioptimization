module F267 (VV235V , VV266V , VV267V); 
input VV235V , VV266V;
output VV267V;
or f0 (VV267V , VV235V , VV266V);
endmodule