module F391 (VV387V , VV390V , VV391V); 
input VV387V , VV390V;
output VV391V;
or f0 (VV391V , VV387V , VV390V);
endmodule