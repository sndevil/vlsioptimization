module F282 (VV278V , VV281V , VV282V); 
input VV278V , VV281V;
output VV282V;
and f0 (VV282V , VV278V , VV281V);
endmodule