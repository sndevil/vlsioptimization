module F68 (VV64V , VV67V , VV68V); 
input VV64V , VV67V;
output VV68V;
or f0 (VV68V , VV64V , VV67V);
endmodule