module F23 (a , d , VV23V); 
input a , d;
output VV23V;
or f0 (VV23V , a , d);
endmodule