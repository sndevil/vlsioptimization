module F395 (VV331V , VV394V , VV395V); 
input VV331V , VV394V;
output VV395V;
or f0 (VV395V , VV331V , VV394V);
endmodule