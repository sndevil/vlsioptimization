module F257 (VV253V , VV256V , VV257V); 
input VV253V , VV256V;
output VV257V;
and f0 (VV257V , VV253V , VV256V);
endmodule