module F20 (e , b , VV20V); 
input e , b;
output VV20V;
and f0 (VV20V , e , b);
endmodule