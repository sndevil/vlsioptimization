module F277 (e , a , VV277V); 
input e , a;
output VV277V;
xor f0 (VV277V , e , a);
endmodule