module F37 (VV35V , VV36V , VV37V); 
input VV35V , VV36V;
output VV37V;
and f0 (VV37V , VV35V , VV36V);
endmodule