module F335 (b , e , VV335V); 
input b , e;
output VV335V;
or f0 (VV335V , b , e);
endmodule