module F66 (d , b , VV66V); 
input d , b;
output VV66V;
or f0 (VV66V , d , b);
endmodule