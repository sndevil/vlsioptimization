module F147 (VV145V , VV146V , VV147V); 
input VV145V , VV146V;
output VV147V;
and f0 (VV147V , VV145V , VV146V);
endmodule