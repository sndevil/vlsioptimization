module F24 (c , d , VV24V); 
input c , d;
output VV24V;
or f0 (VV24V , c , d);
endmodule