module F308 (c , b , VV308V); 
input c , b;
output VV308V;
xor f0 (VV308V , c , b);
endmodule