module F222 (VV220V , VV221V , VV222V); 
input VV220V , VV221V;
output VV222V;
and f0 (VV222V , VV220V , VV221V);
endmodule