module F298 (VV290V , VV297V , VV298V); 
input VV290V , VV297V;
output VV298V;
or f0 (VV298V , VV290V , VV297V);
endmodule