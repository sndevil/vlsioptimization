module F129 (a , d , VV129V); 
input a , d;
output VV129V;
or f0 (VV129V , a , d);
endmodule