module F4 (VV2V , VV3V , VV4V); 
input VV2V , VV3V;
output VV4V;
xor f0 (VV4V , VV2V , VV3V);
endmodule