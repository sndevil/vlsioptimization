module F370 (c , b , VV370V); 
input c , b;
output VV370V;
or f0 (VV370V , c , b);
endmodule