module F210 (VV208V , VV209V , VV210V); 
input VV208V , VV209V;
output VV210V;
and f0 (VV210V , VV208V , VV209V);
endmodule