module F273 (c , b , VV273V); 
input c , b;
output VV273V;
xor f0 (VV273V , c , b);
endmodule