module F388 (e , b , VV388V); 
input e , b;
output VV388V;
xor f0 (VV388V , e , b);
endmodule