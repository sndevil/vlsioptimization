module F97 (VV95V , VV96V , VV97V); 
input VV95V , VV96V;
output VV97V;
or f0 (VV97V , VV95V , VV96V);
endmodule