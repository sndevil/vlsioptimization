module F12 (c , a , VV12V); 
input c , a;
output VV12V;
or f0 (VV12V , c , a);
endmodule