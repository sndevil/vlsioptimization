module F (