module F314 (VV306V , VV313V , VV314V); 
input VV306V , VV313V;
output VV314V;
or f0 (VV314V , VV306V , VV313V);
endmodule