module F135 (b , a , VV135V); 
input b , a;
output VV135V;
or f0 (VV135V , b , a);
endmodule