module F16 (c , e , VV16V); 
input c , e;
output VV16V;
or f0 (VV16V , c , e);
endmodule