module F144 (VV142V' , VV143V , VV144V); 
input VV142V' , VV143V;
output VV144V;
and f0 (VV144V , VV142V' , VV143V);
endmodule