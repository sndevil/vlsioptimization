module F189 (a , c , VV189V); 
input a , c;
output VV189V;
and f0 (VV189V , a , c);
endmodule