module F33 (a , e , VV33V); 
input a , e;
output VV33V;
or f0 (VV33V , a , e);
endmodule