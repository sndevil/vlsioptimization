module F359 (VV357V , VV358V , VV359V); 
input VV357V , VV358V;
output VV359V;
xor f0 (VV359V , VV357V , VV358V);
endmodule