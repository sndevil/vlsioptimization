module F287 (a , e , VV287V); 
input a , e;
output VV287V;
and f0 (VV287V , a , e);
endmodule