module F68 (c , e , VV68V); 
input c , e;
output VV68V;
or f0 (VV68V , c , e);
endmodule