module F217 (VV215V , VV216V , VV217V); 
input VV215V , VV216V;
output VV217V;
or f0 (VV217V , VV215V , VV216V);
endmodule